//module reg_file(input logic Clk, LD, Reset,
//					 input logic[15:0] D,
//					 input logic[2:0] SR2, SR1_M, DR_M,
//					 output logic[15:0] SR1_O, SR2_O);
//always_ff @ (posedge Clk)
//begin
//	if(Reset)
//		SR1_O<=16'h0000;
//		SR2_O<=16'h0000;
//	else 
//		SR1_O<=16h'0000;
//		SR2_O<=16'h0000;
//
//end
//endmodule
